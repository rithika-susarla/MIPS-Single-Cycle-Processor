`timescale 1ns / 1ps

module barrel_shifter(

    );
endmodule
